module mux3 #(parameter WIDTH=8) (a, b, c, select, out);
  // select | out
  // 00 | a
  // 01 | b
  // 02 | c
endmodule
