module simon1 (clock, reset, in, out);
// in:
// R 00
// G 01
// B 10
// Y 11

// out:
// X 00
// 0 01
// 1 10
endmodule
